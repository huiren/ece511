module predict #(parameter WEIGHT_NUM = 33)
(
	input [31:0] ghr,
	input [WEIGHT_NUM*9-1:0] p,
	output logic pred
);

logic [8:0] sum;

always_comb
begin
	sum = p[8:0] // biased
		+ (ghr[0] ? p[17:9] : (~(p[17:9]) + 9'd1))
		+ (ghr[1] ? p[26:18] : (~(p[26:18]) + 9'd1))
		+ (ghr[2] ? p[35:27] : (~(p[35:27]) + 9'd1))
		+ (ghr[3] ? p[44:36] : (~(p[44:36]) + 9'd1))
		+ (ghr[4] ? p[53:45] : (~(p[53:45]) + 9'd1))
		+ (ghr[5] ? p[62:54] : (~(p[62:54]) + 9'd1))
		+ (ghr[6] ? p[71:63] : (~(p[71:63]) + 9'd1))
		+ (ghr[7] ? p[80:72] : (~(p[80:72]) + 9'd1))
		+ (ghr[8] ? p[89:81] : (~(p[89:81]) + 9'd1))
		+ (ghr[9] ? p[98:90] : (~(p[98:90]) + 9'd1))
		+ (ghr[10] ? p[107:99] : (~(p[107:99]) + 9'd1))
		+ (ghr[11] ? p[116:108] : (~(p[116:108]) + 9'd1))
		+ (ghr[12] ? p[125:117] : (~(p[125:117]) + 9'd1))
		+ (ghr[13] ? p[134:126] : (~(p[134:126]) + 9'd1))
		+ (ghr[14] ? p[143:135] : (~(p[143:135]) + 9'd1))
		+ (ghr[15] ? p[152:144] : (~(p[152:144]) + 9'd1))
		+ (ghr[16] ? p[161:153] : (~(p[161:153]) + 9'd1))
		+ (ghr[17] ? p[170:162] : (~(p[170:162]) + 9'd1))
		+ (ghr[18] ? p[179:171] : (~(p[179:171]) + 9'd1))
		+ (ghr[19] ? p[188:180] : (~(p[188:180]) + 9'd1))
		+ (ghr[20] ? p[197:189] : (~(p[197:189]) + 9'd1))
		+ (ghr[21] ? p[206:198] : (~(p[206:198]) + 9'd1))
		+ (ghr[22] ? p[215:207] : (~(p[215:207]) + 9'd1))
		+ (ghr[23] ? p[224:216] : (~(p[224:216]) + 9'd1))
		+ (ghr[24] ? p[233:225] : (~(p[233:225]) + 9'd1))
		+ (ghr[25] ? p[242:234] : (~(p[242:234]) + 9'd1))
		+ (ghr[26] ? p[251:243] : (~(p[251:243]) + 9'd1))
		+ (ghr[27] ? p[260:252] : (~(p[260:252]) + 9'd1))
		+ (ghr[28] ? p[269:261] : (~(p[269:261]) + 9'd1))
		+ (ghr[29] ? p[278:270] : (~(p[278:270]) + 9'd1))
		+ (ghr[30] ? p[287:279] : (~(p[287:279]) + 9'd1))
		+ (ghr[31] ? p[296:288] : (~(p[296:288]) + 9'd1));
end

assign pred = sum[8];

endmodule : predict
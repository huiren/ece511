module predict #(parameter WEIGHT_NUM = 17)
(
	input [15:0] ghr,
	input [WEIGHT_NUM*8-1:0] p,
	output logic pred
);

logic [7:0] sum;

always_comb
begin
	sum = p[7:0] // biased
		+ (ghr[0] ? p[15:8] : (~(p[15:8]) + 8'd1))
		+ (ghr[1] ? p[23:16] : (~(p[23:16]) + 8'd1))
		+ (ghr[2] ? p[31:24] : (~(p[31:24]) + 8'd1))
		+ (ghr[3] ? p[39:32] : (~(p[39:32]) + 8'd1))
		+ (ghr[4] ? p[47:40] : (~(p[47:40]) + 8'd1))
		+ (ghr[5] ? p[55:48] : (~(p[55:48]) + 8'd1))
		+ (ghr[6] ? p[63:56] : (~(p[63:56]) + 8'd1))
		+ (ghr[7] ? p[71:64] : (~(p[71:64]) + 8'd1))
		+ (ghr[8] ? p[79:72] : (~(p[79:72]) + 8'd1))
		+ (ghr[9] ? p[87:80] : (~(p[87:80]) + 8'd1))
		+ (ghr[10] ? p[95:88] : (~(p[95:88]) + 8'd1))
		+ (ghr[11] ? p[103:96] : (~(p[103:96]) + 8'd1))
		+ (ghr[12] ? p[111:104] : (~(p[111:104]) + 8'd1))
		+ (ghr[13] ? p[119:112] : (~(p[119:112]) + 8'd1))
		+ (ghr[14] ? p[127:120] : (~(p[127:120]) + 8'd1))
		+ (ghr[15] ? p[135:128] : (~(p[135:128]) + 8'd1));
end

assign pred = sum[7];

endmodule : predict
